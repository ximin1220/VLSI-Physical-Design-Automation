/users/course/2025F/VLSIPDA202510/g314553017/HW1/lef/asap7sc7p5t_28_SL_4x_220121a.lef