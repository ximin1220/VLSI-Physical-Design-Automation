/users/course/2025F/VLSIPDA202510/g314553017/HW1/lef/asap7_tech_4x_201209.lef